Are the calls are non blocking
Time        Var
0           a
5           c
10          b
20          d
