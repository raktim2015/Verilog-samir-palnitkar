As the calls are blocking, 
Time        Var
0           a
10          b
15          c
35          d
